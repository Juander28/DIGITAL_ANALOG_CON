magic
tech sky130A
magscale 1 2
timestamp 1762817646
<< nwell >>
rect 28843 37257 30254 37910
rect 29538 36300 30138 36621
rect 29818 25824 30161 26124
rect 30078 18684 30142 18748
rect 30470 18354 30534 18418
rect 37366 16469 40608 16482
rect 32722 16402 32786 16466
rect 35144 16206 35208 16270
rect 36079 15443 40608 16469
rect 37366 14402 40608 15443
rect 42736 14402 45918 16482
rect 37599 12066 39240 13092
<< psubdiff >>
rect 28760 20409 31212 20443
<< locali >>
rect 35291 16537 35463 16571
rect 37687 16537 38163 16571
rect 38129 16463 38163 16537
rect 38129 16429 38283 16463
rect 37023 15480 37193 15514
rect 38378 15438 38450 15510
<< viali >>
rect 32737 16417 32771 16451
<< metal1 >>
rect 20776 44364 20856 44392
rect 51654 44364 51714 44370
rect 20776 44304 20784 44364
rect 20844 44304 51654 44364
rect 20776 44290 20856 44304
rect 51654 44298 51714 44304
rect 45568 44130 45652 44140
rect 21784 44070 45581 44130
rect 45641 44070 45652 44130
rect 21784 43636 21844 44070
rect 45568 44058 45652 44070
rect 33945 43826 34005 43832
rect 25626 43766 25632 43826
rect 25692 43766 33945 43826
rect 33945 43760 34005 43766
rect 21776 43626 21854 43636
rect 21776 43566 21784 43626
rect 21844 43566 21854 43626
rect 21776 43556 21854 43566
rect 39170 42784 39242 42790
rect 22248 42724 22254 42784
rect 22314 42724 39176 42784
rect 39236 42724 39242 42784
rect 39170 42718 39242 42724
rect 34356 42408 34428 42414
rect 25202 42348 25208 42408
rect 25268 42348 34362 42408
rect 34422 42348 34428 42408
rect 34356 42342 34428 42348
rect 30078 41538 30142 41544
rect 29467 41486 29473 41538
rect 29525 41526 29531 41538
rect 30078 41526 30084 41538
rect 29525 41498 30084 41526
rect 29525 41486 29531 41498
rect 30078 41486 30084 41498
rect 30136 41486 30142 41538
rect 30078 41480 30142 41486
rect 30269 41194 30333 41200
rect 29302 41142 29308 41194
rect 29360 41182 29366 41194
rect 30269 41182 30275 41194
rect 29360 41154 30275 41182
rect 29360 41142 29366 41154
rect 30269 41142 30275 41154
rect 30327 41142 30333 41194
rect 30269 41136 30333 41142
rect 30476 40992 30528 40998
rect 28955 40940 28961 40992
rect 29013 40980 29019 40992
rect 29013 40952 30476 40980
rect 29013 40940 29019 40952
rect 30476 40934 30528 40940
rect 30078 31301 30141 31307
rect 29473 31249 29479 31301
rect 29531 31289 29537 31301
rect 30078 31289 30084 31301
rect 29531 31261 30084 31289
rect 29531 31249 29537 31261
rect 30078 31249 30084 31261
rect 30136 31249 30141 31301
rect 30078 31243 30141 31249
rect 29309 31121 29361 31127
rect 30269 31121 30332 31127
rect 30269 31109 30275 31121
rect 29361 31081 30275 31109
rect 29309 31063 29361 31069
rect 30269 31069 30275 31081
rect 30327 31069 30332 31121
rect 30269 31063 30332 31069
rect 30470 30946 30534 30952
rect 28955 30894 28961 30946
rect 29013 30934 29019 30946
rect 30470 30934 30476 30946
rect 29013 30906 30476 30934
rect 29013 30894 29019 30906
rect 30470 30894 30476 30906
rect 30528 30894 30534 30946
rect 30470 30888 30534 30894
rect 35164 21276 35224 21282
rect 35164 21210 35224 21216
rect 35164 20848 35224 20854
rect 35164 20782 35224 20788
rect 30078 18742 30142 18748
rect 29468 18690 29474 18742
rect 29526 18730 29532 18742
rect 30078 18730 30084 18742
rect 29526 18702 30084 18730
rect 29526 18690 29532 18702
rect 30078 18690 30084 18702
rect 30136 18690 30142 18742
rect 30078 18684 30142 18690
rect 29312 18576 29364 18582
rect 30275 18576 30327 18582
rect 29364 18536 30275 18564
rect 29312 18518 29364 18524
rect 30275 18518 30327 18524
rect 28966 18412 29018 18418
rect 30470 18412 30534 18418
rect 30470 18400 30476 18412
rect 29018 18372 30476 18400
rect 28966 18354 29018 18360
rect 30470 18360 30476 18372
rect 30528 18360 30534 18412
rect 30470 18354 30534 18360
rect 30856 17088 50842 17160
rect 35164 16716 35224 16722
rect 35164 16650 35224 16656
rect 38376 16580 38452 16592
rect 38376 16528 38388 16580
rect 38440 16528 38452 16580
rect 38376 16516 38452 16528
rect 43288 16520 43294 16572
rect 43346 16520 43352 16572
rect 37730 16472 37794 16478
rect 32722 16460 32786 16466
rect 32722 16408 32728 16460
rect 32780 16408 32786 16460
rect 32722 16402 32786 16408
rect 33382 16460 33434 16466
rect 37730 16420 37736 16472
rect 37788 16420 37794 16472
rect 37730 16414 37794 16420
rect 33382 16402 33434 16408
rect 28521 15400 30911 15534
rect 37025 15470 37194 15522
rect 38378 15504 38450 15510
rect 38378 15444 38384 15504
rect 38444 15444 38450 15504
rect 38378 15438 38450 15444
rect 26602 11056 26608 11236
rect 26788 11056 26794 11236
<< via1 >>
rect 20784 44304 20844 44364
rect 51654 44304 51714 44364
rect 45581 44070 45641 44130
rect 25632 43766 25692 43826
rect 33945 43766 34005 43826
rect 21784 43566 21844 43626
rect 22254 42724 22314 42784
rect 39176 42724 39236 42784
rect 25208 42348 25268 42408
rect 34362 42348 34422 42408
rect 29473 41486 29525 41538
rect 30084 41486 30136 41538
rect 29308 41142 29360 41194
rect 30275 41142 30327 41194
rect 28961 40940 29013 40992
rect 30476 40940 30528 40992
rect 29479 31249 29531 31301
rect 30084 31249 30136 31301
rect 29309 31069 29361 31121
rect 30275 31069 30327 31121
rect 28961 30894 29013 30946
rect 30476 30894 30528 30946
rect 35164 21216 35224 21276
rect 35164 20788 35224 20848
rect 29474 18690 29526 18742
rect 30084 18690 30136 18742
rect 29312 18524 29364 18576
rect 30275 18524 30327 18576
rect 28966 18360 29018 18412
rect 30476 18360 30528 18412
rect 35164 16656 35224 16716
rect 38388 16528 38440 16580
rect 43294 16520 43346 16572
rect 32728 16451 32780 16460
rect 32728 16417 32737 16451
rect 32737 16417 32771 16451
rect 32771 16417 32780 16451
rect 32728 16408 32780 16417
rect 33382 16408 33434 16460
rect 37736 16420 37788 16472
rect 35150 16212 35202 16264
rect 38384 15444 38444 15504
rect 26608 11056 26788 11236
<< metal2 >>
rect 25129 44498 25204 44509
rect 25129 44438 25140 44498
rect 25196 44438 26704 44498
rect 25129 44431 25204 44438
rect 20784 44364 20844 44370
rect 20784 44295 20844 44304
rect 24353 44228 24362 44288
rect 24418 44228 25691 44288
rect 25631 43832 25691 44228
rect 26338 44282 26398 44291
rect 26338 43944 26398 44226
rect 25631 43826 25692 43832
rect 25631 43766 25632 43826
rect 25631 43760 25692 43766
rect 21776 43626 21854 43636
rect 21776 43566 21784 43626
rect 21844 43566 21854 43626
rect 21776 43556 21854 43566
rect 22254 42784 22314 42790
rect 22249 42724 22254 42784
rect 22314 42724 22323 42784
rect 22254 42718 22314 42724
rect 25208 42408 25268 42414
rect 25208 42339 25268 42348
rect 25631 42156 25691 43760
rect 26338 42164 26398 43770
rect 26644 42816 26704 44438
rect 51656 44364 51712 44371
rect 51648 44304 51654 44364
rect 51714 44304 51720 44364
rect 51656 44297 51712 44304
rect 29307 44166 29363 44175
rect 29307 44101 29363 44110
rect 45568 44130 45652 44140
rect 28965 43902 29021 43911
rect 28965 43837 29021 43846
rect 26622 42798 26704 42816
rect 26622 42742 26636 42798
rect 26692 42742 26704 42798
rect 26622 42726 26704 42742
rect 25624 42100 25633 42156
rect 25689 42100 25698 42156
rect 26331 42108 26340 42164
rect 26396 42108 26405 42164
rect 26338 42106 26398 42108
rect 25631 42098 25691 42100
rect 26644 41918 26704 42726
rect 26637 41862 26646 41918
rect 26702 41862 26711 41918
rect 28979 41886 29007 43837
rect 26644 41860 26704 41862
rect 29321 41856 29349 44101
rect 45568 44070 45581 44130
rect 45641 44070 45652 44130
rect 45568 44058 45652 44070
rect 33939 43824 33945 43826
rect 34005 43824 34011 43826
rect 33938 43768 33945 43824
rect 34005 43768 34012 43824
rect 33939 43766 33945 43768
rect 34005 43766 34011 43768
rect 39170 42784 39242 42790
rect 39170 42782 39176 42784
rect 39236 42782 39242 42784
rect 39169 42726 39176 42782
rect 39236 42726 39243 42782
rect 39170 42724 39176 42726
rect 39236 42724 39242 42726
rect 39170 42718 39242 42724
rect 34356 42408 34428 42414
rect 34356 42406 34362 42408
rect 34422 42406 34428 42408
rect 29477 42366 29533 42375
rect 34355 42350 34362 42406
rect 34422 42350 34429 42406
rect 34356 42348 34362 42350
rect 34422 42348 34428 42350
rect 34356 42342 34428 42348
rect 29477 42301 29533 42310
rect 29740 42324 29796 42333
rect 29491 41842 29519 42301
rect 29740 42259 29796 42268
rect 29754 41932 29782 42259
rect 29762 41661 29882 41689
rect 29473 41538 29525 41544
rect 29473 41480 29525 41486
rect 30078 41538 30142 41544
rect 30078 41486 30084 41538
rect 30136 41486 30142 41538
rect 30078 41480 30142 41486
rect 29308 41194 29360 41200
rect 29308 41136 29360 41142
rect 30269 41194 30333 41200
rect 30269 41142 30275 41194
rect 30327 41142 30333 41194
rect 30269 41136 30333 41142
rect 28961 40992 29013 40998
rect 30470 40940 30476 40992
rect 30528 40940 30534 40992
rect 28961 40934 29013 40940
rect 29771 31406 29882 31434
rect 29479 31301 29531 31307
rect 29479 31243 29531 31249
rect 30078 31301 30141 31307
rect 30078 31249 30084 31301
rect 30136 31249 30141 31301
rect 30078 31243 30141 31249
rect 30269 31121 30332 31127
rect 29303 31069 29309 31121
rect 29361 31069 29367 31121
rect 30269 31069 30275 31121
rect 30327 31069 30332 31121
rect 30269 31063 30332 31069
rect 28961 30946 29013 30952
rect 28961 30888 29013 30894
rect 30470 30946 30534 30952
rect 30470 30894 30476 30946
rect 30528 30894 30534 30946
rect 30470 30888 30534 30894
rect 35166 21276 35222 21283
rect 35158 21216 35164 21276
rect 35224 21216 35230 21276
rect 35166 21209 35222 21216
rect 35158 20846 35164 20848
rect 35224 20846 35230 20848
rect 35157 20790 35164 20846
rect 35224 20790 35231 20846
rect 35158 20788 35164 20790
rect 35224 20788 35230 20790
rect 29759 19332 29882 19360
rect 29474 18742 29526 18748
rect 29474 18684 29526 18690
rect 30078 18742 30142 18748
rect 30078 18690 30084 18742
rect 30136 18690 30142 18742
rect 30078 18684 30142 18690
rect 29306 18524 29312 18576
rect 29364 18524 29370 18576
rect 30269 18524 30275 18576
rect 30327 18524 30333 18576
rect 30470 18412 30534 18418
rect 28960 18360 28966 18412
rect 29018 18360 29024 18412
rect 30470 18360 30476 18412
rect 30528 18360 30534 18412
rect 30470 18354 30534 18360
rect 35158 16714 35164 16716
rect 35224 16714 35230 16716
rect 35157 16658 35164 16714
rect 35224 16658 35231 16714
rect 35158 16656 35164 16658
rect 35224 16656 35230 16658
rect 38376 16582 38452 16592
rect 38376 16526 38386 16582
rect 38442 16526 38452 16582
rect 38376 16516 38452 16526
rect 43294 16572 43346 16578
rect 43294 16514 43346 16520
rect 37730 16472 37794 16478
rect 37730 16469 37736 16472
rect 32722 16460 32786 16466
rect 32722 16408 32728 16460
rect 32780 16451 32786 16460
rect 33376 16451 33382 16460
rect 32780 16417 33382 16451
rect 32780 16408 32786 16417
rect 33376 16408 33382 16417
rect 33434 16408 33440 16460
rect 35153 16423 37736 16469
rect 32722 16402 32786 16408
rect 35153 16270 35199 16423
rect 37730 16420 37736 16423
rect 37788 16469 37794 16472
rect 43297 16469 43343 16514
rect 37788 16423 43343 16469
rect 37788 16420 37794 16423
rect 37730 16414 37794 16420
rect 35144 16264 35208 16270
rect 35144 16212 35150 16264
rect 35202 16212 35208 16264
rect 35144 16206 35208 16212
rect 38378 15504 38450 15510
rect 38378 15502 38384 15504
rect 38444 15502 38450 15504
rect 38377 15446 38384 15502
rect 38444 15446 38451 15502
rect 38378 15444 38384 15446
rect 38444 15444 38450 15446
rect 38378 15438 38450 15444
rect 26608 11236 26788 11242
rect 26608 9388 26788 11056
rect 26498 9208 26788 9388
rect 26498 8059 26678 9208
rect 26494 7889 26503 8059
rect 26673 7889 26682 8059
rect 26498 7884 26678 7889
<< via2 >>
rect 25140 44438 25196 44498
rect 20784 44304 20844 44360
rect 24362 44228 24418 44288
rect 26338 44226 26398 44282
rect 21784 43566 21844 43626
rect 22258 42724 22314 42784
rect 25208 42348 25268 42404
rect 51656 44306 51712 44362
rect 29307 44110 29363 44166
rect 28965 43846 29021 43902
rect 26636 42742 26692 42798
rect 25633 42100 25689 42156
rect 26340 42108 26396 42164
rect 26646 41862 26702 41918
rect 45583 44072 45639 44128
rect 33947 43768 34003 43824
rect 39178 42726 39234 42782
rect 29477 42310 29533 42366
rect 34364 42350 34420 42406
rect 29740 42268 29796 42324
rect 35166 21218 35222 21274
rect 35166 20790 35222 20846
rect 35166 16658 35222 16714
rect 38386 16580 38442 16582
rect 38386 16528 38388 16580
rect 38388 16528 38440 16580
rect 38440 16528 38442 16580
rect 38386 16526 38442 16528
rect 38386 15446 38442 15502
rect 26503 7889 26673 8059
<< metal3 >>
rect 25107 44503 25220 44525
rect 25107 44439 25135 44503
rect 25201 44439 25220 44503
rect 25107 44438 25140 44439
rect 25196 44438 25220 44439
rect 25107 44408 25220 44438
rect 20760 44363 20866 44392
rect 20760 44299 20779 44363
rect 20849 44299 20866 44363
rect 51651 44362 51717 44367
rect 51651 44306 51656 44362
rect 51712 44306 51717 44362
rect 51651 44301 51717 44306
rect 20760 44280 20866 44299
rect 24000 44226 24006 44290
rect 24070 44288 24076 44290
rect 24357 44288 24423 44293
rect 24070 44228 24362 44288
rect 24418 44228 24423 44288
rect 24070 44226 24076 44228
rect 24357 44223 24423 44228
rect 24904 44286 24968 44292
rect 26330 44284 26336 44290
rect 24968 44226 26336 44284
rect 26400 44226 26406 44290
rect 24968 44224 26403 44226
rect 24904 44216 24968 44222
rect 26333 44221 26403 44224
rect 21794 44204 21858 44210
rect 29730 44192 29736 44256
rect 29800 44192 29806 44256
rect 21794 44134 21858 44140
rect 20792 44006 20856 44012
rect 7922 43944 20792 44004
rect 7922 41918 7982 43944
rect 20792 43936 20856 43942
rect 21796 43636 21856 44134
rect 26810 44106 26816 44170
rect 26880 44168 26886 44170
rect 29302 44168 29368 44171
rect 26880 44166 29368 44168
rect 26880 44110 29307 44166
rect 29363 44110 29368 44166
rect 26880 44108 29368 44110
rect 26880 44106 26886 44108
rect 29302 44105 29368 44108
rect 25212 44060 25276 44066
rect 22268 44038 22332 44044
rect 29467 43996 29473 44060
rect 29537 43996 29543 44060
rect 25212 43990 25276 43996
rect 22268 43968 22332 43974
rect 21776 43626 21856 43636
rect 21776 43624 21784 43626
rect 13995 43566 21784 43624
rect 21844 43566 21856 43626
rect 13995 43564 21856 43566
rect 13995 41848 14055 43564
rect 21776 43556 21854 43564
rect 22270 42789 22330 43968
rect 22253 42784 22330 42789
rect 22253 42758 22258 42784
rect 20400 42724 22258 42758
rect 22314 42724 22330 42784
rect 20400 42698 22330 42724
rect 20400 41856 20460 42698
rect 25214 42409 25274 43990
rect 25994 43842 26000 43906
rect 26064 43904 26070 43906
rect 28960 43904 29026 43907
rect 26064 43902 29026 43904
rect 26064 43846 28965 43902
rect 29021 43846 29026 43902
rect 26064 43844 29026 43846
rect 26064 43842 26070 43844
rect 28960 43841 29026 43844
rect 25720 43634 25784 43640
rect 25714 43572 25720 43632
rect 25784 43572 26852 43632
rect 25720 43564 25784 43570
rect 26606 42802 26732 42822
rect 26606 42738 26632 42802
rect 26696 42738 26732 42802
rect 26606 42716 26732 42738
rect 25203 42404 25274 42409
rect 25203 42348 25208 42404
rect 25268 42348 25274 42404
rect 26792 42366 26852 43572
rect 29475 42371 29535 43996
rect 29472 42366 29538 42371
rect 25203 42343 25274 42348
rect 25214 41880 25274 42343
rect 26784 42302 26790 42366
rect 26854 42302 26860 42366
rect 29472 42310 29477 42366
rect 29533 42310 29538 42366
rect 29738 42329 29798 44192
rect 45568 44128 45652 44140
rect 45568 44072 45583 44128
rect 45639 44072 45652 44128
rect 45568 44058 45652 44072
rect 33942 43824 34008 43829
rect 33942 43768 33947 43824
rect 34003 43768 34008 43824
rect 33942 43763 34008 43768
rect 33230 43540 33236 43604
rect 33300 43540 33306 43604
rect 30018 42738 30024 42802
rect 30088 42800 30094 42802
rect 30088 42740 32992 42800
rect 30088 42738 30094 42740
rect 30044 42582 30108 42588
rect 32782 42582 32846 42588
rect 30108 42520 32782 42580
rect 30044 42512 30108 42518
rect 32782 42512 32846 42518
rect 29472 42305 29538 42310
rect 29735 42324 29801 42329
rect 29735 42268 29740 42324
rect 29796 42268 29801 42324
rect 29735 42263 29801 42268
rect 26335 42164 26401 42169
rect 25628 42156 25694 42161
rect 25628 42100 25633 42156
rect 25689 42100 25694 42156
rect 26335 42108 26340 42164
rect 26396 42108 26401 42164
rect 26335 42103 26401 42108
rect 25628 42095 25694 42100
rect 25631 41904 25691 42095
rect 26338 41872 26398 42103
rect 26641 41918 26707 41923
rect 26641 41862 26646 41918
rect 26702 41862 26707 41918
rect 26641 41857 26707 41862
rect 32932 41854 32992 42740
rect 33238 41854 33298 43540
rect 33945 41876 34005 43763
rect 38087 43001 38093 43199
rect 38291 43001 38297 43199
rect 39170 42782 39242 42790
rect 39170 42726 39178 42782
rect 39234 42726 39242 42782
rect 39170 42718 39242 42726
rect 34356 42406 34428 42414
rect 34356 42350 34364 42406
rect 34420 42350 34428 42406
rect 34356 42342 34428 42350
rect 34362 41900 34422 42342
rect 39176 41850 39236 42718
rect 45581 41828 45641 44058
rect 51654 42046 51714 44301
rect 35161 21274 35227 21279
rect 35161 21218 35166 21274
rect 35222 21218 35227 21274
rect 35161 21213 35227 21218
rect 35164 20851 35224 21213
rect 35161 20846 35227 20851
rect 35161 20790 35166 20846
rect 35222 20790 35227 20846
rect 35161 20785 35227 20790
rect 30661 18784 30725 18790
rect 30661 18714 30725 18720
rect 35164 16719 35224 20785
rect 35161 16714 35227 16719
rect 35161 16658 35166 16714
rect 35222 16658 35227 16714
rect 35161 16653 35227 16658
rect 38376 16582 38452 16592
rect 38376 16526 38386 16582
rect 38442 16526 38452 16582
rect 38376 16516 38452 16526
rect 38384 15510 38444 16516
rect 38378 15502 38450 15510
rect 38378 15446 38386 15502
rect 38442 15446 38450 15502
rect 38378 15438 38450 15446
rect 26498 8059 26678 8064
rect 26498 7889 26503 8059
rect 26673 7889 26678 8059
rect 26498 6969 26678 7889
rect 26498 6791 26499 6969
rect 26677 6791 26678 6969
rect 26498 6790 26678 6791
rect 26499 6785 26677 6790
rect 537 5526 935 5531
rect 536 5525 56328 5526
rect 536 5127 537 5525
rect 935 5467 56328 5525
rect 935 5455 28154 5467
rect 935 5429 24768 5455
rect 935 5425 16450 5429
rect 935 5413 12158 5425
rect 935 5373 7460 5413
rect 935 5175 4074 5373
rect 4272 5215 7460 5373
rect 7658 5401 12158 5413
rect 7658 5215 9464 5401
rect 4272 5203 9464 5215
rect 9662 5371 12158 5401
rect 9662 5203 10154 5371
rect 4272 5175 10154 5203
rect 935 5173 10154 5175
rect 10352 5227 12158 5371
rect 12356 5395 16450 5425
rect 12356 5227 15544 5395
rect 10352 5197 15544 5227
rect 15742 5231 16450 5395
rect 16648 5409 24768 5429
rect 16648 5401 21840 5409
rect 16648 5231 18454 5401
rect 15742 5203 18454 5231
rect 18652 5211 21840 5401
rect 22038 5395 24768 5409
rect 22038 5211 22764 5395
rect 18652 5203 22764 5211
rect 15742 5197 22764 5203
rect 22962 5257 24768 5395
rect 24966 5269 28154 5455
rect 28352 5463 56328 5467
rect 28352 5461 43894 5463
rect 28352 5447 37598 5461
rect 28352 5377 36674 5447
rect 28352 5269 31284 5377
rect 24966 5257 31284 5269
rect 22962 5197 31284 5257
rect 10352 5179 31284 5197
rect 31482 5249 36674 5377
rect 36872 5263 37598 5447
rect 37796 5455 43894 5461
rect 37796 5263 40984 5455
rect 36872 5257 40984 5263
rect 41182 5407 43894 5455
rect 41182 5257 42988 5407
rect 36872 5249 42988 5257
rect 31482 5209 42988 5249
rect 43186 5265 43894 5407
rect 44092 5461 56328 5463
rect 44092 5441 55364 5461
rect 44092 5265 47280 5441
rect 43186 5243 47280 5265
rect 47478 5433 55364 5441
rect 47478 5243 49284 5433
rect 43186 5235 49284 5243
rect 49482 5405 55364 5433
rect 49482 5349 51978 5405
rect 49482 5235 49974 5349
rect 43186 5209 49974 5235
rect 31482 5179 49974 5209
rect 10352 5173 49974 5179
rect 935 5151 49974 5173
rect 50172 5207 51978 5349
rect 52176 5263 55364 5405
rect 55562 5263 56328 5461
rect 52176 5207 56328 5263
rect 50172 5151 56328 5207
rect 935 5127 56328 5151
rect 536 5126 56328 5127
rect 537 5121 935 5126
<< via3 >>
rect 25135 44498 25201 44503
rect 25135 44439 25140 44498
rect 25140 44439 25196 44498
rect 25196 44439 25201 44498
rect 20779 44360 20849 44363
rect 20779 44304 20784 44360
rect 20784 44304 20844 44360
rect 20844 44304 20849 44360
rect 20779 44299 20849 44304
rect 24006 44226 24070 44290
rect 24904 44222 24968 44286
rect 26336 44282 26400 44290
rect 26336 44226 26338 44282
rect 26338 44226 26398 44282
rect 26398 44226 26400 44282
rect 21794 44140 21858 44204
rect 29736 44192 29800 44256
rect 20792 43942 20856 44006
rect 26816 44106 26880 44170
rect 22268 43974 22332 44038
rect 25212 43996 25276 44060
rect 29473 43996 29537 44060
rect 26000 43842 26064 43906
rect 25720 43570 25784 43634
rect 26632 42798 26696 42802
rect 26632 42742 26636 42798
rect 26636 42742 26692 42798
rect 26692 42742 26696 42798
rect 26632 42738 26696 42742
rect 26790 42302 26854 42366
rect 33236 43540 33300 43604
rect 30024 42738 30088 42802
rect 30044 42518 30108 42582
rect 32782 42518 32846 42582
rect 38093 43001 38291 43199
rect 30661 18720 30725 18784
rect 26499 6791 26677 6969
rect 537 5127 935 5525
rect 4074 5175 4272 5373
rect 7460 5215 7658 5413
rect 9464 5203 9662 5401
rect 10154 5173 10352 5371
rect 12158 5227 12356 5425
rect 15544 5197 15742 5395
rect 16450 5231 16648 5429
rect 18454 5203 18652 5401
rect 21840 5211 22038 5409
rect 22764 5197 22962 5395
rect 24768 5257 24966 5455
rect 28154 5269 28352 5467
rect 31284 5179 31482 5377
rect 36674 5249 36872 5447
rect 37598 5263 37796 5461
rect 40984 5257 41182 5455
rect 42988 5209 43186 5407
rect 43894 5265 44092 5463
rect 47280 5243 47478 5441
rect 49284 5235 49482 5433
rect 49974 5151 50172 5349
rect 51978 5207 52176 5405
rect 55364 5263 55562 5461
<< metal4 >>
rect 200 5526 600 44152
rect 1612 43444 2012 44152
rect 6134 43444 6194 45152
rect 6686 43444 6746 45152
rect 7238 43444 7298 45152
rect 7790 43444 7850 45152
rect 8342 43444 8402 45152
rect 8894 43444 8954 45152
rect 9446 43444 9506 45152
rect 9998 43444 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44392 21650 45152
rect 20776 44363 21650 44392
rect 20776 44299 20779 44363
rect 20849 44332 21650 44363
rect 20849 44299 20856 44332
rect 20776 44290 20856 44299
rect 20794 44007 20854 44290
rect 21793 44204 21859 44205
rect 21793 44140 21794 44204
rect 21858 44202 21859 44204
rect 22142 44202 22202 45152
rect 21858 44142 22202 44202
rect 21858 44140 21859 44142
rect 21793 44139 21859 44140
rect 22267 44038 22333 44039
rect 20791 44006 20857 44007
rect 20791 43942 20792 44006
rect 20856 43942 20857 44006
rect 22267 43974 22268 44038
rect 22332 44036 22333 44038
rect 22694 44036 22754 45152
rect 23246 44058 23306 45152
rect 23798 44288 23858 45152
rect 24005 44290 24071 44291
rect 24005 44288 24006 44290
rect 23798 44228 24006 44288
rect 24005 44226 24006 44228
rect 24070 44226 24071 44290
rect 24005 44225 24071 44226
rect 24350 44284 24410 45152
rect 24902 44501 24962 45152
rect 25134 44503 25202 44504
rect 25134 44501 25135 44503
rect 24902 44441 25135 44501
rect 25134 44439 25135 44441
rect 25201 44439 25202 44503
rect 25134 44438 25202 44439
rect 24903 44286 24969 44287
rect 24903 44284 24904 44286
rect 24350 44224 24904 44284
rect 24903 44222 24904 44224
rect 24968 44222 24969 44286
rect 24903 44221 24969 44222
rect 25211 44060 25277 44061
rect 25211 44058 25212 44060
rect 22332 43976 22754 44036
rect 23244 43998 25212 44058
rect 25211 43996 25212 43998
rect 25276 43996 25277 44060
rect 25211 43995 25277 43996
rect 22332 43974 22333 43976
rect 22267 43973 22333 43974
rect 20791 43941 20857 43942
rect 25454 43632 25514 45152
rect 26006 43982 26066 45152
rect 26335 44290 26401 44291
rect 26335 44226 26336 44290
rect 26400 44226 26401 44290
rect 26335 44225 26401 44226
rect 26002 43907 26066 43982
rect 25999 43906 26066 43907
rect 25999 43842 26000 43906
rect 26064 43878 26066 43906
rect 26064 43842 26065 43878
rect 25999 43841 26065 43842
rect 25719 43634 25785 43635
rect 25719 43632 25720 43634
rect 25454 43572 25720 43632
rect 25719 43570 25720 43572
rect 25784 43570 25785 43634
rect 25719 43569 25785 43570
rect 26338 43602 26398 44225
rect 26558 44168 26618 45152
rect 26815 44170 26881 44171
rect 26815 44168 26816 44170
rect 26558 44110 26816 44168
rect 26562 44108 26816 44110
rect 26815 44106 26816 44108
rect 26880 44106 26881 44170
rect 26815 44105 26881 44106
rect 27110 44058 27170 45152
rect 27662 44254 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 29735 44256 29801 44257
rect 29735 44254 29736 44256
rect 27662 44194 29736 44254
rect 29735 44192 29736 44194
rect 29800 44192 29801 44256
rect 29735 44191 29801 44192
rect 29472 44060 29538 44061
rect 29472 44058 29473 44060
rect 27110 43998 29473 44058
rect 29472 43996 29473 43998
rect 29537 43996 29538 44060
rect 29472 43995 29538 43996
rect 33235 43604 33301 43605
rect 33235 43602 33236 43604
rect 26338 43542 33236 43602
rect 33235 43540 33236 43542
rect 33300 43540 33301 43604
rect 33235 43539 33301 43540
rect 1612 43199 55674 43444
rect 1612 43044 38093 43199
rect 200 5525 936 5526
rect 200 5127 537 5525
rect 935 5127 936 5525
rect 200 5126 936 5127
rect 200 1000 600 5126
rect 1612 1000 2012 43044
rect 4621 39474 4821 43044
rect 8454 39494 8654 43044
rect 14224 39520 14424 43044
rect 15543 43042 15743 43044
rect 15543 40686 15743 41618
rect 16449 40730 16649 41620
rect 18069 39488 18269 43044
rect 21344 39532 21544 43044
rect 26048 39744 26248 43044
rect 26622 42802 26704 42816
rect 26622 42738 26632 42802
rect 26696 42800 26704 42802
rect 30023 42802 30089 42803
rect 30023 42800 30024 42802
rect 26696 42740 30024 42800
rect 26696 42738 26704 42740
rect 26622 42726 26704 42738
rect 30023 42738 30024 42740
rect 30088 42738 30089 42802
rect 30023 42737 30089 42738
rect 30043 42582 30109 42583
rect 30043 42580 30044 42582
rect 27386 42520 30044 42580
rect 26789 42366 26855 42367
rect 26789 42302 26790 42366
rect 26854 42302 26855 42366
rect 26789 42301 26855 42302
rect 26792 42210 26852 42301
rect 27386 42210 27446 42520
rect 30043 42518 30044 42520
rect 30108 42518 30109 42582
rect 30043 42517 30109 42518
rect 26792 42150 27446 42210
rect 26792 41850 26852 42150
rect 31730 39518 31930 43044
rect 32781 42582 32847 42583
rect 32781 42518 32782 42582
rect 32846 42518 32847 42582
rect 32781 42517 32847 42518
rect 32784 41910 32844 42517
rect 33388 39678 33588 43044
rect 38092 43001 38093 43044
rect 38291 43044 55674 43199
rect 38291 43001 38292 43044
rect 38092 39518 38292 43001
rect 41367 39488 41567 43044
rect 45212 39486 45412 43044
rect 50982 39512 51182 43044
rect 54815 39496 55015 43044
rect 30660 18784 30726 18785
rect 30660 18720 30661 18784
rect 30725 18720 30726 18784
rect 30660 18719 30726 18720
rect 4073 5373 4273 13910
rect 4073 5175 4074 5373
rect 4272 5175 4273 5373
rect 7459 5413 7659 13034
rect 7459 5215 7460 5413
rect 7658 5215 7659 5413
rect 7459 5214 7659 5215
rect 9463 5401 9663 13800
rect 9463 5203 9464 5401
rect 9662 5203 9663 5401
rect 9463 5202 9663 5203
rect 10153 5371 10353 14538
rect 4073 5174 4273 5175
rect 10153 5173 10154 5371
rect 10352 5173 10353 5371
rect 12157 5425 12357 14516
rect 12157 5227 12158 5425
rect 12356 5227 12357 5425
rect 12157 5226 12357 5227
rect 15543 5395 15743 12868
rect 15543 5197 15544 5395
rect 15742 5197 15743 5395
rect 16449 5429 16649 12888
rect 16449 5231 16450 5429
rect 16648 5231 16649 5429
rect 16449 5230 16649 5231
rect 18453 5401 18653 12606
rect 18453 5203 18454 5401
rect 18652 5203 18653 5401
rect 21839 5409 22039 12694
rect 21839 5211 21840 5409
rect 22038 5211 22039 5409
rect 21839 5210 22039 5211
rect 22763 5395 22963 12646
rect 18453 5202 18653 5203
rect 15543 5196 15743 5197
rect 22763 5197 22764 5395
rect 22962 5197 22963 5395
rect 24767 5455 24967 12688
rect 24767 5257 24768 5455
rect 24966 5257 24967 5455
rect 24767 5256 24967 5257
rect 26498 6969 26678 6970
rect 26498 6791 26499 6969
rect 26677 6791 26678 6969
rect 22763 5196 22963 5197
rect 10153 5172 10353 5173
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 6791
rect 28153 5467 28353 12708
rect 28153 5269 28154 5467
rect 28352 5269 28353 5467
rect 28153 5268 28353 5269
rect 30663 1830 30723 18719
rect 31283 5377 31483 18192
rect 31730 15496 31930 17614
rect 33388 15496 33588 17494
rect 31283 5179 31284 5377
rect 31482 5179 31483 5377
rect 34669 5192 34869 18164
rect 36673 5447 36873 18216
rect 36673 5249 36674 5447
rect 36872 5249 36873 5447
rect 37597 5461 37797 18460
rect 37597 5263 37598 5461
rect 37796 5263 37797 5461
rect 37597 5262 37797 5263
rect 40983 5455 41183 18402
rect 36673 5248 36873 5249
rect 40983 5257 40984 5455
rect 41182 5257 41183 5455
rect 31283 5178 31483 5179
rect 40983 5136 41183 5257
rect 42987 5407 43187 18366
rect 42987 5209 42988 5407
rect 43186 5209 43187 5407
rect 43893 5463 44093 18352
rect 43893 5265 43894 5463
rect 44092 5265 44093 5463
rect 43893 5264 44093 5265
rect 47279 5441 47479 18408
rect 47279 5243 47280 5441
rect 47478 5243 47479 5441
rect 47279 5234 47479 5243
rect 49283 5433 49483 18210
rect 49283 5235 49284 5433
rect 49482 5235 49483 5433
rect 49283 5234 49483 5235
rect 49973 5349 50173 18240
rect 42987 5150 43187 5209
rect 49973 5151 49974 5349
rect 50172 5151 50173 5349
rect 51977 5405 52177 18330
rect 51977 5207 51978 5405
rect 52176 5207 52177 5405
rect 55363 5461 55563 18272
rect 55363 5263 55364 5461
rect 55562 5263 55563 5461
rect 55363 5262 55563 5263
rect 51977 5206 52177 5207
rect 49973 5150 50173 5151
rect 30362 1770 30723 1830
rect 30362 0 30542 1770
use BASIC_SQRT  BASIC_SQRT_0 ~/Documents/GERMAN/magic/SQRT
timestamp 1762682500
transform 1 0 29542 0 -1 18337
box 4782 -3330 15196 2911
use BASIC_SQRT  BASIC_SQRT_1
timestamp 1762682500
transform -1 0 58440 0 -1 18337
box 4782 -3330 15196 2911
use BASIC_SQRT  BASIC_SQRT_2
timestamp 1762682500
transform 1 0 23854 0 1 12532
box 4782 -3330 15196 2911
use BASIC_SQRT  BASIC_SQRT_3
timestamp 1762682500
transform 1 0 23680 0 -1 14957
box 4782 -3330 15196 2911
use BDW5  BDW5_0 ~/Documents/GERMAN/magic/BDW
timestamp 1762796168
transform 1 0 29768 0 1 38815
box 42 -21674 26310 3346
use BDW6  BDW6_0 ~/Documents/GERMAN/magic/BDW
timestamp 1762795706
transform -1 0 29868 0 1 38815
box 29 -26619 26308 3346
use CON_IV_phvt_nn  CON_IV_phvt_nn_0 ~/Documents/GERMAN/magic/CON_IV_HVT
timestamp 1760947506
transform 1 0 25889 0 -1 18315
box 4928 1212 11216 2872
use CON_IV_phvt_nn  CON_IV_phvt_nn_1
timestamp 1760947506
transform -1 0 56058 0 1 12556
box 4928 1212 11216 2872
use CON_IV_phvt_nn  CON_IV_phvt_nn_2
timestamp 1760947506
transform -1 0 33768 0 1 9338
box 4928 1212 11216 2872
use CON_IV_phvt_nn  CON_IV_phvt_nn_3
timestamp 1760947506
transform -1 0 49744 0 1 12556
box 4928 1212 11216 2872
use CON_IV_phvt_nn  CON_IV_phvt_nn_4
timestamp 1760947506
transform -1 0 49430 0 -1 14938
box 4928 1212 11216 2872
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 1612 1000 2012 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
